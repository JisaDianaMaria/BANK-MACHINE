library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
entity afisare_contalegere is
	port(	  
	      enable:in  std_logic; 
		   clk:in  std_logic:='0';	
	      c1: in  std_logic_vector(1 downto 0); 
	      catod:  out std_logic_vector(6 downto 0);	
		   an:  out std_logic_vector(3 downto 0));
end entity;
 
architecture bcdsegm of afisare_contalegere is
signal cifra: std_logic_vector(1 downto 0);
signal counter: std_logic_vector(1 downto 0):="00";
begin		
  										 
	process(cifra)
	begin
		case cifra is
				when "00" =>  catod<="0000001"; --0
				when "01" =>  catod<="1001111"; --1
				when "10" =>  catod<="0010010"; --2
				when "11" =>  catod<="0000110"; --3
			    when others => catod<="1111111";
			end case;
	end process;	
	process(clk,enable)
	begin
		if(clk='1' and clk'event and enable='1') then 
		        case counter is 
				    when "00"=>  cifra<="00";
					 when "01"=>  cifra<="00";
				    when "10"=>  cifra<="00"; 
			       when others => cifra<=c1;
			 end case;	   
		
        end if;
	     
	end process;
  process(clk)
       begin
            if(clk='1' and clk'event) then
               counter<=counter +1;
            end if;     
       end process;
	 process(counter)
       begin
            case counter  is
                when "00" => an<="0111";
                when "01" => an<="1011";
                when "10" => an<="1101";
                when others => an<="1110";
             
            end case;
       end process;   
end architecture;